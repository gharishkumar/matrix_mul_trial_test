module adder16(a, b, clk, sum);
    input [15:0] a, b;
    input clk;
    output reg [15:0] sum;

    always @(posedge clk) begin
        sum <= a + b;
    end
endmodule